* RC Filter Testbench
* -------------------
.control
  pre_osdi rc_filter.osdi    ; load your Verilog-A model
  run                        ; run the simulation

  set filetype=ascii         ; make the raw file readable text
  write rc_filter.raw all    ; save all simulation data

  plot v(in) v(out)          ; plot both signals in the GUI
  hardcopy rc_filter.eps v(in) v(out)


  quit
.endc

Vin in 0 SIN(0 1 1k)

.model myrc rc_filter R=1000 C=1e-6
N1 in out myrc

Rload out 0 1e6

.tran 1us 5ms
.end
